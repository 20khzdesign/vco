volt to octave 

.include ../../../spice/AD8519.cir
.include ../../../spice/LM741.cir


.SUBCKT OPAMP1	     1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* GAIN BW PRODUCT = 10MHZ
* DC GAIN (100K) AND POLE 1 (100HZ)
EGAIN	3 0	1 2	100K
RP1	3	4	1K
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS

vin key 0 DC 1V

r1   key   3    5k
r2   3     in   10k

X1   0   3   in   OPAMP1
