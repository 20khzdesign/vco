OPINV.CIR - OPAMP INVERTING AMPLIFIER
*
VS	1	0	AC	1	SIN(0V	1VPEAK	10KHZ)
*
R1	1	2	5K
R2	2	4	10K
XOP	0 2	4	OPAMP1	
*
* OPAMP MACRO MODEL, SINGLE-POLE 
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1	     1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* GAIN BW PRODUCT = 10MHZ
* DC GAIN (100K) AND POLE 1 (100HZ)
EGAIN	3 0	1 2	100K
RP1	3	4	1K
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS
*
* ANALYSIS 
.AC 	DEC 	5 1K 10MEG
.TRAN 	0.005MS  0.2MS
* VIEW RESULTS
.PRINT	AC 	VM(1) VM(4)
.PLOT	AC 	VM(1) VM(4)
.PRINT	TRAN 	V(1) V(4)
.PLOT	TRAN 	V(1) V(4)
.PROBE
.END
